`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/07 14:57:40
// Design Name: 
// Module Name: Master
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Master(
    // Global Signals
    input logic clk,
    input logic reset,
    // Button Interface
    input logic run_stop,
    input logic clear,
    // SPI Interface
    output logic o_SCLK,
    output logic o_MOSI,
    output logic o_SS_N, 
    input logic i_MISO     // �̹� ������Ʈ������ FND Controll�� �����̴ٺ���, ��������� ����.

    );

    // Internal Signals
    logic [7:0] tx_data;
    logic start;
    logic ss_n;
    logic tx_ready;
    logic done;

    SPI_Master U_SPI_Master (
        .clk(clk),
        .reset(reset),
        .start(start),
        .tx_data(tx_data),
        .tx_ready(tx_ready),
        .done(done),
        .SCLK(o_SCLK),
        .MOSI(o_MOSI),
        .MISO(i_MISO)
    );

    // SS_N�� UpCounter���� ���� ����
    assign o_SS_N = ss_n;

    UpCounter U_UpCounter (
        .clk(clk),
        .reset(reset),
        .run_stop(run_stop),
        .clear(clear),
        .tx_ready(tx_ready),
        .done(done),
        .tx_data(tx_data),
        .start(start),
        .ss_n(ss_n)
    );
endmodule





module UpCounter(
    // Global Signals
    input logic clk,
    input logic reset,
    // Input Signals (Buttons)
    input logic run_stop,    // ī��Ʈ ����/���� ���
    input logic clear,       // ī���� �ʱ�ȭ
    // Input Signals (From SPI Master)
    input logic tx_ready,    // SPI Master�� ���� �غ� �Ϸ� (IDLE ����)
    input logic done,        // SPI Master�� ���� �Ϸ� (8bit ���� ��)
    // Output Signals (To SPI Master)
    output logic [7:0] tx_data,   // ������ 8bit ������ (0~255)
    output logic start,           // SPI ���� ���� ��ȣ
    output logic ss_n             // Slave Select ��ȣ (Active Low)
    );

    // ========================================
    // ��ǥ ����:
    // 1. run_stop ��ư: ī��Ʈ ����/���� ���
    // 2. clear ��ư: ī���� 0���� �ʱ�ȭ
    // 3. 8��Ʈ ī���� (0~255 �ݺ�)
    // 4. ���� �ֱ�� ī��Ʈ ���� �� SPI ����
    // 5. tx_ready Ȯ�� �� start ��ȣ �߻� (�浹 ����)
    // 6. done ��ȣ�� ���� �Ϸ� Ȯ��
    // ========================================

    typedef enum logic [3:0] {
        IDLE,
        RUN,
        STOP,
        CLEAR_SEND,        // Clear �� ��� 0 ����
        WAIT_TX_READY,
        SEND_HIGH_BYTE,
        WAIT_HIGH_DONE,
        SEND_LOW_BYTE,
        WAIT_LOW_DONE
    } state_t;

    state_t c_state, n_state;

    // Registers
    logic [13:0] counter_reg, counter_next;      // 14��Ʈ ī���� (0~9999)
    logic [31:0] clk_count_reg, clk_count_next;  // �ֱ� ī��Ʈ��
    logic start_reg, start_next;                  // SPI ���� ��ȣ
    logic ss_n_reg, ss_n_next;                   // Slave Select ��ȣ
    logic return_to_idle_reg, return_to_idle_next; // ���� �Ϸ� �� IDLE�� ���ư��� ����

    // ========================================
    // State Register
    // ========================================
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            c_state <= IDLE;
            counter_reg <= 14'd0;
            clk_count_reg <= 32'd0;
            start_reg <= 1'b0;
            ss_n_reg <= 1'b1;  // SS_N = High (��Ȱ��)
            return_to_idle_reg <= 1'b0;
        end else begin
            c_state <= n_state;
            counter_reg <= counter_next;
            clk_count_reg <= clk_count_next;
            start_reg <= start_next;
            ss_n_reg <= ss_n_next;
            return_to_idle_reg <= return_to_idle_next;
        end
    end

    // ========================================
    // Next State Logic + Output Logic
    // ========================================
    always_comb begin
        // �⺻�� ���� (Latch ����)
        n_state = c_state;
        counter_next = counter_reg;
        clk_count_next = clk_count_reg;
        start_next = 1'b0;
        ss_n_next = 1'b1;  // �⺻��: SS_N = High (��Ȱ��)
        return_to_idle_next = return_to_idle_reg;
        
        case(c_state)
            IDLE: begin
                // �ʱ� ����: ī���� ����
                counter_next = 14'd0;
                clk_count_next = 32'd0;
                start_next = 1'b0;
                
                if (clear) begin
                    n_state = CLEAR_SEND;  // Clear �� ��� 0 ����
                end else if (run_stop) begin
                    n_state = RUN;
                end else begin
                    n_state = IDLE;
                end
            end

            RUN: begin
                // ī���� ��: ���� �ֱ⸶�� ����
                if (clear) begin
                    // Clear ��ư: ��� �ʱ�ȭ �� 0 ����
                    counter_next = 14'd0;
                    clk_count_next = 32'd0;
                    n_state = CLEAR_SEND;
                end else if (run_stop) begin
                    // Run/Stop ��ư: ���� �� �����ϰ� ����
                    clk_count_next = 32'd0;
                    n_state = STOP;
                end else begin
                    // ���� �ֱ� üũ (��: 0.01�ʸ��� ���� = 1,000,000 Ŭ��)
                    if (clk_count_reg >= 32'd9_999_999) begin
                        clk_count_next = 32'd0;
                        // 14��Ʈ ī����: 0~9999 ��ȯ
                        if (counter_reg >= 14'd9999) begin
                            counter_next = 14'd0;
                        end else begin
                            counter_next = counter_reg + 1'b1;
                        end
                        n_state = WAIT_TX_READY;  // SPI ���� �غ�
                    end else begin
                        clk_count_next = clk_count_reg + 1'b1;
                        n_state = RUN;
                    end
                end
            end

            STOP: begin
                // ���� ����: ī���� �� ����
                counter_next = counter_reg;
                clk_count_next = 32'd0;
                start_next = 1'b0;
                
                if (clear) begin
                    counter_next = 14'd0;
                    n_state = CLEAR_SEND;  // Clear �� ��� 0 ����
                end else if (run_stop) begin
                    n_state = RUN;
                end else begin
                    n_state = STOP;
                end
            end

            CLEAR_SEND: begin
                // *** Clear ��ư �� ��� 0 ���� ***
                // counter_reg�� �̹� 0���� ������
                counter_next = 14'd0;
                clk_count_next = 32'd0;
                start_next = 1'b0;
                ss_n_next = 1'b1;  // ���� ��Ȱ��
                return_to_idle_next = 1'b1;  // ���� �Ϸ� �� IDLE�� ����
                
                // SPI Master�� �غ�Ǹ� ��� 0 ����
                if (tx_ready) begin
                    n_state = SEND_HIGH_BYTE;  // 0 �� ���� ����
                end else begin
                    n_state = CLEAR_SEND;  // �غ�� ������ ���
                end
            end

            WAIT_TX_READY: begin
                // *** SPI Master�� �غ�� ������ ��� ***
                // tx_ready=1�̸� SPI Master�� IDLE ���� (���� ����)
                start_next = 1'b0;
                ss_n_next = 1'b1;  // ���� ��Ȱ��
                return_to_idle_next = 1'b0;  // ���� ī�����̹Ƿ� RUN���� ����
                
                if (tx_ready) begin
                    n_state = SEND_HIGH_BYTE;  // ���� ����Ʈ ���� ����
                end else begin
                    n_state = WAIT_TX_READY;  // ��� ���
                end
            end

            SEND_HIGH_BYTE: begin
                // *** ���� ����Ʈ ���� ���� ***
                start_next = 1'b1;  // start �޽� (1Ŭ��)
                ss_n_next = 1'b0;   // SS_N = Low (Slave Ȱ��ȭ)
                n_state = WAIT_HIGH_DONE;
            end

            WAIT_HIGH_DONE: begin
                // *** ���� ����Ʈ ���� �Ϸ� ��� ***
                start_next = 1'b0;  // start ��ȣ ����
                ss_n_next = 1'b0;   // SS_N = Low ���� (���� ���� ��)
                
                if (done) begin
                    n_state = SEND_LOW_BYTE;  // ���� ����Ʈ �������� �̵�
                end else begin
                    n_state = WAIT_HIGH_DONE;  // ���� �Ϸ���� ���
                end
            end

            SEND_LOW_BYTE: begin
                // *** ���� ����Ʈ ���� ���� ***
                start_next = 1'b1;  // start �޽� (1Ŭ��)
                ss_n_next = 1'b0;   // SS_N = Low ����
                n_state = WAIT_LOW_DONE;
            end

            WAIT_LOW_DONE: begin
                // *** ���� ����Ʈ ���� �Ϸ� ��� ***
                start_next = 1'b0;  // start ��ȣ ����
                ss_n_next = 1'b0;   // SS_N = Low ����
                
                if (done) begin
                    ss_n_next = 1'b1;  // ��� ���� �Ϸ� �� SS_N = High (��Ȱ��ȭ)
                    // ���� �Ϸ� �� ���ư� ���� ����
                    if (return_to_idle_reg) begin
                        n_state = IDLE;  // Clear���� �� ��� IDLE��
                    end else begin
                        n_state = RUN;   // ���� ī���ÿ��� �� ��� RUN����
                    end
                end else begin
                    n_state = WAIT_LOW_DONE;  // ���� �Ϸ���� ���
                end
            end

            default: begin
                n_state = IDLE;
                counter_next = 14'd0;
                clk_count_next = 32'd0;
                start_next = 1'b0;
                ss_n_next = 1'b1;  // �⺻��: ��Ȱ��
                return_to_idle_next = 1'b0;
            end
        endcase
    end

    // ========================================
    // ��� �Ҵ�
    // ========================================
    // 2-byte ����: ���� ����Ʈ�� ���� ����Ʈ ����
    // counter_reg: 0~9999 �� High:��������Ʈ(counter/100), Low:��������Ʈ(counter%100)
    logic [7:0] high_byte, low_byte;
    assign high_byte = counter_reg / 100;    // ����: 0~99 (100�� �ڸ�)
    assign low_byte = counter_reg % 100;     // ����: 0~99 (1�� �ڸ�)
    
    // ���� ���¿� ���� ������ ����Ʈ ����
    assign tx_data = (c_state == SEND_HIGH_BYTE || c_state == WAIT_HIGH_DONE) ? high_byte : low_byte;
    assign start = start_reg;
    assign ss_n = ss_n_reg;             // SS_N ��ȣ ���

endmodule


module SPI_Master (
    // Global Signals
    input logic clk,
    input logic reset,
    // Internal Signals
    input logic start,
    input logic [7:0] tx_data,
    output logic [7:0] rx_data,
    output logic tx_ready,
    output logic done,
    // External SPI Signals
    output logic SCLK,
    output logic MOSI,
    input logic MISO
    // SS_N�� UpCounter���� ���� ����
);


    // ���� ���迡����, SCLK�� ���ֱ⸦ CPO(SCLK=0), ������ �� �ֱ⸦ CP1(SCLK=1)�� �����ϰ�,
    // �� State���� MOSI, MISO ��ȣ�� ó���ϴ� ������� ����.
    typedef enum {
        IDLE,
        CP0,
        CP1
    } state_t;

    state_t c_state, n_state;

    logic [7:0] tx_data_reg, tx_data_next;          // To prevent Latch
    logic [7:0] rx_data_reg, rx_data_next;          // To prevent Latch

    logic [5:0] sclk_count_reg, sclk_count_next;    // To prevent Latch
    logic [2:0] bit_count_reg, bit_count_next;        // To prevent Latch


    // State Register
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            c_state <= IDLE;
            tx_data_reg <= 8'b0;
            rx_data_reg <= 8'b0;
            sclk_count_reg <= 6'b0;
            bit_count_reg <= 3'b0;
        end else begin
            c_state <= n_state;
            tx_data_reg <= tx_data_next;
            rx_data_reg <= rx_data_next;
            sclk_count_reg <= sclk_count_next;
            bit_count_reg <= bit_count_next;
        end
    end


    // Next State Logic(Combinational) + Output Logic(Combinational)
    always_comb begin
        n_state = c_state;  // �⺻�� ����
        tx_data_next = tx_data_reg;  // �⺻�� ����
        rx_data_next = rx_data_reg;  // �⺻�� ����
        sclk_count_next = sclk_count_reg;  // �⺻�� ����
        bit_count_next = bit_count_reg;  // �⺻�� ����
        tx_ready = 1'b0;  // �⺻�� ����
        done = 1'b0;  // �⺻�� ����
        SCLK = 1'b0;  // CPOL = 0����, �⺻�� ����
        case (c_state)
            IDLE: begin
                    done = 1'b0;          // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                    tx_ready = 1'b1;      // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                    sclk_count_next = 0;
                    bit_count_next = 0;
                if (start) begin
                    n_state = CP0;
                    tx_data_next = tx_data;  //TX data latching
                end else begin
                    n_state = IDLE;
                end
            end
            CP0: begin
                SCLK = 0; // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                if (sclk_count_reg == 49) begin    // Rising Edge
                    rx_data_next = {rx_data_reg[6:0], MISO};  // MSB first ����
                    sclk_count_next = 0;
                    n_state = CP1;
                end else begin
                    sclk_count_next = sclk_count_reg + 1;
                    n_state = CP0;
                end
            end
            CP1: begin
                SCLK = 1; // Output Port ��ȣ�̹Ƿ�, registerȭ ���� �ʾƵ� ��.
                if (sclk_count_reg == 49) begin
                    sclk_count_next = 0;
                    if (bit_count_reg == 7) begin   // Falling Edge
                        bit_count_next = 0;
                        done = 1;
                        n_state = IDLE;
                    end else begin
                        bit_count_next = bit_count_reg + 1;
                        tx_data_next = {tx_data_reg[6:0], 1'b0};  // MSB first ����
                        n_state = CP0;
                    end
                end else begin
                    sclk_count_next = sclk_count_reg + 1;
                    n_state = CP1;
                end
            end
        endcase
    end

    // ��, tx_data, bit_count, sclk_count���� ��ȣ���� ��������ȭ �ߴ°�?
    // => Latch ���� ����.
    // => Combinational logic���� ��ȣ�� ���� ���¸� ������ ��,
    //    �ش� ��ȣ���� ��������ȭ �Ǿ� ���� ������, ��ȣ�� ���� ���¸� �����ϱ� ���� Latch�� ������ �� ����.
    //    �̴� ����ġ ���� ������ �ʷ��� �� ����.
    // ������ ���� �ش� ��ȣ�� Module�� output ��Ʈ���, ��������ȭ ���� �ʾƵ� ��.
    // => Module�� output ��Ʈ�� �⺻������ Combinational logic���� ���� �Ҵ�ޱ� ������,
    //    Latch�� ������ ������ ����. 
    //
    // ��, ����� internal signal���� combinational logic�ӿ��� �� ���� �ٲ�� �ȴٸ�
    // �ش� signal���� ��������ȭ �ؾ���. (LATCH ���� ����)
    // �ݸ鿡, ����� output ��Ʈ���� ��������ȭ ���� �ʾƵ� ��.

    assign MOSI = tx_data_reg[7];  // MSB first ����
    assign rx_data = rx_data_reg;  // ���� ���� ������
endmodule
