`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/07 15:00:51
// Design Name: 
// Module Name: Slave
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Slave(
    // Global Signals
    input logic clk,
    input logic reset,
    // SPI Interface (��� FPGA�� Master�κ��� ������ ��ȣ)
    input logic i_SCLK,
    input logic i_MOSI,
    input logic i_SS_N, 
    output logic o_MISO,
    // Fnd Interface
    output logic [6:0] fnd_data,
    output logic [3:0] fnd_com
    );

    // Internal Signals
    logic [7:0] w_rx_data;    // SPI Slave�� ������ ������
    logic w_done;              // SPI ���� �Ϸ� ��ȣ
    logic [13:0] w_fnd_data;   // FND ǥ�ÿ� 14bit ������


    SPI_Slave U_SPI_Slave (
        .clk(clk),
        .reset(reset),
        .i_SCLK(i_SCLK),
        .i_MOSI(i_MOSI),
        .i_SS_N(i_SS_N),
        .o_MISO(o_MISO),
        .rx_data(w_rx_data),
        .done(w_done)
    );

    ControlUnit U_ControlUnit (
        .clk(clk),
        .reset(reset),
        .rx_data(w_rx_data),
        .done(w_done),
        .fnd_data(w_fnd_data)
    );

    fnd_controller U_Fnd_controller (
        .clk(clk),
        .rst(reset),
        .i_fnd_data(w_fnd_data),
        .o_fnd_data(fnd_data),
        .fnd_com(fnd_com)
    );

endmodule


module SPI_Slave(
    // Global Signals
    input logic clk,          // System clock (FPGA ���� Ŭ�� - 100MHz)
    input logic reset,
    // SPI Interface (�ܺ� Master�κ��� ������ ��ȣ��)
    input logic i_SCLK,       // Master�κ��� �޴� SPI Clock (���� Ŭ��, ��: 1MHz)
    input logic i_MOSI,       // Master�κ��� �޴� ������ (Master Out Slave In)
    input logic i_SS_N,       // Slave Select (Active Low - 0�� �� Ȱ��ȭ)
    output logic o_MISO,      // Master���� ������ ������ (Master In Slave Out, ���� �̻��)
    // Control Unit Interface
    output logic [7:0] rx_data,  // ���� �Ϸ�� 8bit ������
    output logic done            // ���� �Ϸ� ��ȣ (1Ŭ�� �޽�)
    );

    // ========================================
    // Slave�� �ܺο��� ������ SCLK�� ����ȭ�Ǿ�� ��
    // ������ �ý��� Ŭ��(clk)���� �����ϸ鼭 SCLK�� edge�� �����ϴ� ��� ���
    // ========================================
    
    // SCLK�� SS_N ����ȭ �������� (Metastability ������)
    logic [2:0] sclk_sync;     // 3�ܰ� ����ȭ (CDC - Clock Domain Crossing)
    logic [2:0] ss_n_sync;     // 3�ܰ� ����ȭ
    
    // Edge detection ��ȣ
    logic sclk_rising_edge;    // SCLK�� 0->1 ��ȭ ����
    logic sclk_falling_edge;   // SCLK�� 1->0 ��ȭ ����
    logic ss_n_active;          // SS_N�� Ȱ��ȭ(Low) ��������
    
    // Data registers
    logic [7:0] rx_shift_reg;   // ���� ������ ����Ʈ �������� (��Ʈ���� ��ĭ�� �̵�)
    logic [7:0] tx_shift_reg;   // �۽� ������ ����Ʈ �������� (MISO��, ���� �̻��)
    logic [2:0] bit_counter;     // ��Ʈ ī���� (0~7���� ī��Ʈ)
    logic rx_done;              // ���� ���� �Ϸ� �÷���
    
    
    // ========================================
    // 1�ܰ�: SCLK�� SS_N ����ȭ (Metastability ����)
    // ========================================
    // �ܺο��� ������ �񵿱� ��ȣ�� �ý��� Ŭ���� ����ȭ
    // 3�� �ø��÷����� ����ȭ�Ͽ� �������� ��ȣ ����
    // �ϸ�, Synchronizer��� �Ҹ�
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            sclk_sync <= 3'b000;
            ss_n_sync <= 3'b111;  // SS_N�� �⺻������ High (��Ȱ��)
        end else begin
            // 3��Ʈ ����Ʈ �������ͷ� ����ȭ
            sclk_sync <= {sclk_sync[1:0], i_SCLK};  // [2]�� ���� �������� ��ȣ
            ss_n_sync <= {ss_n_sync[1:0], i_SS_N};
        end
    end
    
    // Edge detection: ���� ��(bit[2])�� ���� ��(bit[1])�� ��
    assign sclk_rising_edge = (sclk_sync[2:1] == 2'b01);   // 0->1 transition
    assign sclk_falling_edge = (sclk_sync[2:1] == 2'b10);  // 1->0 transition
    assign ss_n_active = ~ss_n_sync[2];  // Active Low�̹Ƿ� ���� (0�� �� true)
    
    
    // ========================================
    // 2�ܰ�: SPI Slave ���� ���� (CPOL=0, CPHA=0 ����)
    // ========================================
    // SPI ���: CPOL=0 (Idle ���¿��� SCLK=0), CPHA=0 (ù ��° edge���� ���ø�)
    // ����:
    //   - SCLK Rising Edge (0->1): MOSI �����͸� �о shift register�� ����
    //   - SCLK Falling Edge (1->0): ���� ��Ʈ�� �غ� (MISO ������Ʈ, ���� �̻��)
    //   - 8��Ʈ ���� �Ϸ� �� done ��ȣ �߻�
    
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            rx_shift_reg <= 8'h00;
            tx_shift_reg <= 8'h00;
            bit_counter <= 3'd0;
            rx_done <= 1'b0;
        end 
        else begin
            rx_done <= 1'b0;  // �⺻������ done�� 0 (1Ŭ�� �޽��� ����)
            
            if (!ss_n_active) begin
                // SS_N�� High (��Ȱ��)�̸� �ʱ�ȭ
                // Slave�� ���õ��� ���� ����
                bit_counter <= 3'd0;
                rx_shift_reg <= 8'h00;
                tx_shift_reg <= 8'h00;
            end 
            else begin
                // SS_N�� Low (Ȱ��)�� ���� SPI ��� ����
                
                if (sclk_rising_edge) begin
                    // *** �߿�: SCLK Rising Edge���� MOSI ������ ���ø� ***
                    // MSB First ���: ���� ���� ��Ʈ�� ���� ��Ʈ
                    rx_shift_reg <= {rx_shift_reg[6:0], i_MOSI};  
                    bit_counter <= bit_counter + 1'b1;
                    
                    // 8��Ʈ ��� ���� �Ϸ� (bit 7���� ������ ���� edge���� ī���Ͱ� 0�� ��)
                    if (bit_counter == 3'd7) begin
                        rx_done <= 1'b1;      // ���� �Ϸ� ��ȣ (1Ŭ�� �޽�)
                        bit_counter <= 3'd0;  // ���� ����Ʈ�� ���� ����
                    end
                end
                
                // Falling Edge������ MISO �غ� (���� ������Ʈ������ ��� ����)
                // if (sclk_falling_edge) begin
                //     tx_shift_reg <= {tx_shift_reg[6:0], 1'b0};  // ���� ��Ʈ �غ�
                // end
            end
        end
    end
    
    
    // Output Logic
    assign rx_data = rx_shift_reg;  // ���� ���ŵ� ������ (8��Ʈ �Ϸ� �� ��ȿ)
    assign done = rx_done;           // ���� �Ϸ� ��ȣ (8��Ʈ ���� �Ϸ� �� 1Ŭ�� ���� High)
    
    // MISO�� ���� ������Ʈ���� ������� ���� (�ܹ��� FND Control ����)
    // �ʿ�� tx_shift_reg�� MSB�� ����ϸ� ��
    assign o_MISO = 1'b0;  // �Ǵ� tx_shift_reg[7];
    
endmodule



// ========================================
// Control Unit: SPI�� ���� 2���� 8bit �����͸� �����Ͽ� 0~9999 ǥ��
// ========================================
// 
// *** �ٽ� ���̵��: 2-Byte ���� ***
// - Master�� 0~9999 ���� 2���� 8bit�� �����ؼ� ����
// - ���ڵ� ���: high_byte = value/100, low_byte = value%100
// - ���ڵ� ���: fnd_data = (high_byte �� 100) + low_byte
// 
// ����:
//   1. ù ��° done: rx_data �� high_byte (����: 0~99, 100�� �ڸ�)
//   2. �� ��° done: rx_data �� low_byte (����: 0~99, 1�� �ڸ�)
//   3. fnd_data = high_byte �� 100 + low_byte (0~9999)
//
module ControlUnit(
    input logic clk,
    input logic reset,
    input logic [7:0] rx_data,   // SPI�� ������ 8bit ������ (0~255)
    input logic done,             // SPI ���� �Ϸ� ��ȣ (1Ŭ�� �޽�)
    output logic [13:0] fnd_data  // FND ǥ�ÿ� 14bit ������ (0~9999)
);

    // State machine
    typedef enum logic [1:0] {
        WAIT_HIGH_BYTE,    // ù ��° ����Ʈ (����) ���
        WAIT_LOW_BYTE,     // �� ��° ����Ʈ (����) ���
        UPDATE_DISPLAY     // ���÷��� ������Ʈ
    } state_t;

    state_t c_state, n_state;
    
    // Registers
    logic [7:0] high_byte_reg, high_byte_next;   // ���� ����Ʈ ���� (0~99)
    logic [13:0] fnd_data_reg, fnd_data_next;    // ���� FND ������ (0~9999)

    
    // ========================================
    // State Register
    // ========================================
    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            c_state <= WAIT_HIGH_BYTE;
            high_byte_reg <= 8'd0;
            fnd_data_reg <= 14'd0;
        end else begin
            c_state <= n_state;
            high_byte_reg <= high_byte_next;
            fnd_data_reg <= fnd_data_next;
        end
    end


    // ========================================
    // Next State Logic + Output Logic (Combinational)
    // ========================================
    always_comb begin
        // �⺻�� ���� (Latch ����)
        n_state = c_state;
        high_byte_next = high_byte_reg;
        fnd_data_next = fnd_data_reg;
        
        case(c_state)
            WAIT_HIGH_BYTE: begin
                // ù ��° ����Ʈ (����) ���� ���
                if (done) begin
                    n_state = WAIT_LOW_BYTE;
                    high_byte_next = rx_data;       // ���� ����Ʈ ���� (0~99)
                    fnd_data_next = fnd_data_reg;   // FND ������ ����
                end else begin
                    n_state = WAIT_HIGH_BYTE;
                end
            end

            WAIT_LOW_BYTE: begin
                // �� ��° ����Ʈ (����) ���� ���
                if (done) begin
                    n_state = UPDATE_DISPLAY;
                    
                    // *** �ٽ� ����: (high �� 100) + low ***
                    // high_byte_reg: 0~99 (100�� �ڸ�)
                    // rx_data:       0~99 (1�� �ڸ�)
                    fnd_data_next = (high_byte_reg * 100) + rx_data;
                    
                    // ������ġ: 9999 �ʰ� �� wrapping
                    if (fnd_data_next == 14'd9999) begin
                        fnd_data_next = 14'd0;
                    end
                    
                    high_byte_next = 8'd0;  // ��� �Ϸ�
                end else begin
                    n_state = WAIT_LOW_BYTE;
                end
            end

            UPDATE_DISPLAY: begin
                // ���÷��� ������Ʈ �Ϸ�, ���� ������ ���
                n_state = WAIT_HIGH_BYTE;
            end

            default: begin
                n_state = WAIT_HIGH_BYTE;
                high_byte_next = 8'd0;
                fnd_data_next = 14'd0;
            end
        endcase
    end
    
    // ========================================
    // ���
    // ========================================
    assign fnd_data = fnd_data_reg;

endmodule


// 10000�� couunter
module fnd_controller(
    input [13:0] i_fnd_data,
    input  clk,
    input  rst,
    output [6:0] o_fnd_data,
    output [3:0] fnd_com
    );

    wire [3:0] w_digit_1;
    wire [3:0] w_digit_10;
    wire [3:0] w_digit_100;
    wire [3:0] w_digit_1000;
    wire [3:0] w_bcd;
    wire [1:0] w_digit_sel;

    wire w_1khz;


    digit_spliter U_DS(
        .i_data(i_fnd_data),  
        .digit_1(w_digit_1),
        .digit_10(w_digit_10),
        .digit_100(w_digit_100),
        .digit_1000(w_digit_1000)
    );

    bcd_decoder U_BCD(
        .bcd(w_bcd),
        .fnd_data(o_fnd_data)
    );


    mux_4x1 U_MUX4_1(
        .sel(w_digit_sel),
        .digit_1(w_digit_1),
        .digit_10(w_digit_10),
        .digit_100(w_digit_100),
        .digit_1000(w_digit_1000),
        .bcd_data(w_bcd)
    );
    
    mux_2x4 U_Mux_Fnd_com(
        .sel(w_digit_sel),
        .fnd_com(fnd_com)
    );

    counter_4 U_CNT_4(
        .clk(w_1khz),
        .rst(rst),
        .digit_sel(w_digit_sel)
    );

    clk_div U_CLK_DIV(
        .clk(clk),
        .rst(rst),
        .o_1khz(w_1khz)
    );

endmodule



module digit_spliter(
    input [13:0] i_data,   // 8bit吏쒕?�� sov_e + cov
    
    output [3:0] digit_1,
    output [3:0] digit_10,
    output [3:0] digit_100,
    output [3:0] digit_1000
);

    assign digit_1 = i_data % 10;
    assign digit_10 = i_data/10 % 10;
    assign digit_100 = i_data/100 % 10;
    assign digit_1000 = i_data/1000 % 10;

endmodule


module bcd_decoder(
    input [3:0]bcd,
    output reg [6:0]fnd_data  
);

    always @(bcd) begin
        case(bcd)
            0 : fnd_data =  7'h40;  // 7-bit: 1000000 (segments a,b,c,d,e,f)
            1 : fnd_data =  7'h79;  // 7-bit: 1111001 (segments b,c)
            2 : fnd_data =  7'h24;  // 7-bit: 0100100 (segments a,b,g,e,d)
            3 : fnd_data =  7'h30;  // 7-bit: 0110000 (segments a,b,g,c,d)
            4 : fnd_data =  7'h19;  // 7-bit: 0011001 (segments f,g,b,c)
            5 : fnd_data =  7'h12;  // 7-bit: 0010010 (segments a,f,g,c,d)
            6 : fnd_data =  7'h02;  // 7-bit: 0000010 (segments a,f,g,e,d,c)
            7 : fnd_data =  7'h78;  // 7-bit: 1111000 (segments a,b,c)
            8 : fnd_data =  7'h00;  // 7-bit: 0000000 (all segments)
            9 : fnd_data =  7'h10;  // 7-bit: 0010000 (segments a,b,c,d,f,g)
            default : fnd_data = 7'h7f; // 7-bit: all off
        endcase
    end

endmodule



module mux_4x1(
    input [1:0] sel,
    input [3:0]digit_1,
    input [3:0]digit_10,
    input [3:0]digit_100,        
    input [3:0]digit_1000,    
    output reg [3:0] bcd_data
    );


    always @(*) begin
        case(sel)
            2'b00 : bcd_data = digit_1;
            2'b01 : bcd_data = digit_10;
            2'b10 : bcd_data = digit_100;
            2'b11 : bcd_data = digit_1000;
            default : bcd_data = digit_1;
        endcase
     end    

endmodule

module mux_2x4(
        input [1:0] sel,
        output reg [3:0] fnd_com
    );

    always @(sel) begin
        case(sel)
            2'b00 : fnd_com = 4'b1110;
            2'b01 : fnd_com = 4'b1101;
            2'b10 : fnd_com = 4'b1011;
            2'b11 : fnd_com = 4'b0111;
            default : fnd_com = 4'b1111;
        endcase
    end

    


endmodule

module counter_4(
    input clk,
    input rst,
    output [1:0] digit_sel
    );

    reg [1:0] r_counter;

    assign digit_sel = r_counter;

    always@(posedge clk or posedge rst)begin
        if(rst) begin
            r_counter <= 2'b00;
        end
        else begin
            r_counter <= r_counter + 1'b1;
        end
    end
    
endmodule


module clk_div(
    input clk,
    input rst,
    output reg o_1khz
    );

    reg [16:0]r_counter;

always @(posedge clk or posedge rst)begin
    if(rst) begin
        r_counter <= 0;
        o_1khz <= 0;
    end 
    else begin
    if(r_counter == 100_000-1 ) begin
        r_counter <= 0;
        o_1khz <= 1'b1;
    end
    else begin
        r_counter <= r_counter + 1'b1;
        o_1khz <= 0;
        end
    end
end

endmodule
